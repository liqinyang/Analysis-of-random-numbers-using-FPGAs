module mt_mem(
input clk,
input rst,
input enable,
input [623:0][31:0] in,
output reg [623:0][31:0]out);



always@(posedge clk)
if (rst)begin
	out<={32'd116925273,32'd373236455,32'd538248802,32'd4226154574,32'd1600421663,32'd3144139009,32'd1274635091,32'd4237523457,32'd4127642404,32'd745796080,32'd2898003956,32'd1198755052,32'd996401156,32'd3491702910,32'd1163546293,32'd2185572068,32'd2739416220,32'd864314942,32'd4185309254,32'd1123937393,32'd371107437,32'd1652380747,32'd254886981,32'd2739135905,32'd3160415220,32'd2980581379,32'd2058599240,32'd2605376692,32'd2259549051,32'd939608650,32'd2093376088,32'd559792668,32'd35512535,32'd2601327385,32'd3745016485,32'd1857807303,32'd2134869635,32'd75235680,32'd2192917968,32'd1427007580,32'd68338106,32'd2452128692,32'd3565923316,32'd3846781604,32'd2968478428,32'd3046897033,32'd593715887,32'd3358845388,32'd2112227260,32'd1796963839,32'd3920626153,32'd3165387311,32'd1196168985,32'd2251039304,32'd3710224584,32'd1238643345,32'd4010345846,32'd4089211432,32'd2165639585,32'd2820237500,32'd3477775846,32'd1833692038,32'd182251010,32'd2782204324,32'd3174283928,32'd1339524978,32'd994467513,32'd153529770,32'd755541153,32'd1243290919,32'd1822261341,32'd358193390,32'd1623822350,32'd29887881,32'd562407139,32'd3920910597,32'd3715040333,32'd2773634239,32'd4050094885,32'd2351938991,32'd339011744,32'd1389255297,32'd575756423,32'd1170979324,32'd3039860130,32'd2473777375,32'd1148331655,32'd3672652561,32'd3146108732,32'd1084892922,32'd3920699442,32'd1610171318,32'd841138647,32'd3433623522,32'd3601685135,32'd32037606,32'd2125374725,32'd3712771231,32'd1404047266,32'd3510589272,32'd511679284,32'd4136013972,32'd220376185,32'd4290295859,32'd1481153225,32'd3523379959,32'd4187931679,32'd257453352,32'd1214999983,32'd1824668777,32'd2988544460,32'd3033724173,32'd2593265787,32'd1342921678,32'd1682465785,32'd1273083041,32'd3616954837,32'd2268543712,32'd3381351589,32'd903950702,32'd916922266,32'd2430244594,32'd2534236055,32'd2772611204,32'd4259079565,32'd1212963762,32'd3789435080,32'd439487268,32'd3926825101,32'd2261078634,32'd2844468873,32'd3884997363,32'd3444379103,32'd327684603,32'd2450260579,32'd2514956543,32'd213886228,32'd2527167744,32'd4209506140,32'd1024058911,32'd2035120316,32'd3427511545,32'd1651820702,32'd2796251125,32'd3625937786,32'd1082871720,32'd3242113092,32'd1124291831,32'd2114916962,32'd2801191520,32'd2991889790,32'd1628818384,32'd3105466755,32'd586888764,32'd4102349079,32'd1468131552,32'd841637218,32'd980275996,32'd1207204018,32'd4188936761,32'd4246466163,32'd2747624534,32'd1322770750,32'd678802395,32'd242514037,32'd2604438657,32'd2827490451,32'd357178131,32'd721365878,32'd1894847490,32'd1064389665,32'd4270524229,32'd3279042455,32'd462404995,32'd3207806491,32'd2480850074,32'd2011314805,32'd2932420675,32'd2932285520,32'd3031943234,32'd3411729501,32'd3250223302,32'd3849196601,32'd1040109604,32'd3574242559,32'd719279415,32'd1273496002,32'd2947436871,32'd24441053,32'd3938010494,32'd237854258,32'd3543438633,32'd396985542,32'd284638153,32'd1639223168,32'd4193124145,32'd2140815539,32'd968642107,32'd499920867,32'd2448981354,32'd4198420524,32'd3467616712,32'd1798831929,32'd3173743570,32'd699324101,32'd1641962571,32'd4093330405,32'd3762293788,32'd1153351468,32'd2671701715,32'd1170828427,32'd2317706652,32'd2627897488,32'd2530947598,32'd3741110422,32'd3060733996,32'd1549973222,32'd4226219908,32'd751549633,32'd4126386549,32'd2397606939,32'd1728726693,32'd410962657,32'd3129049475,32'd88291794,32'd3159187032,32'd3718575695,32'd144842260,32'd4070363626,32'd657841564,32'd1225135658,32'd2709796449,32'd746910746,32'd3072795503,32'd605849491,32'd2920887680,32'd1690255681,32'd1995296581,32'd2227353703,32'd2677441952,32'd1499184106,32'd4017453944,32'd526022968,32'd4202067531,32'd2288745211,32'd4277634633,32'd3197046734,32'd3926649337,32'd238724805,32'd1683964498,32'd355877597,32'd1122941824,32'd3306178891,32'd4101820340,32'd10753957,32'd3482428591,32'd3459298550,32'd3346805556,32'd451352804,32'd2395942225,32'd2902374922,32'd1560546623,32'd1484884283,32'd2907371963,32'd1664731394,32'd2787463443,32'd4122051269,32'd3054207519,32'd177954239,32'd635252598,32'd969180562,32'd1601509561,32'd2033930425,32'd660912408,32'd3510695954,32'd4097726412,32'd3876142393,32'd102527300,32'd2545470627,32'd2493306969,32'd2901327722,32'd49780221,32'd2124571119,32'd2213336821,32'd1294126893,32'd2551930098,32'd3110908772,32'd2957657929,32'd3733051177,32'd4233923286,32'd3339845861,32'd2122918776,32'd3444590461,32'd824266620,32'd426751932,32'd93044840,32'd4058078927,32'd3362203896,32'd3467353606,32'd540086248,32'd1123848930,32'd2889497980,32'd2059099269,32'd1780609115,32'd2411256222,32'd539226467,32'd4068324016,32'd1981273229,32'd2683353,32'd3882821767,32'd3742425828,32'd3762283879,32'd3389311029,32'd2534774459,32'd351970715,32'd3779331880,32'd1097832595,32'd636350498,32'd3694851522,32'd2538837125,32'd4148487199,32'd1419478013,32'd3422594099,32'd1879502046,32'd1987859863,32'd3847120877,32'd1187340812,32'd1424193429,32'd2684567658,32'd2356924521,32'd3283991819,32'd818418468,32'd1999436060,32'd1388503581,32'd2448282623,32'd4264711934,32'd3111170404,32'd3209557296,32'd2933843154,32'd4121720519,32'd3029422620,32'd1858551310,32'd1478959417,32'd4294466702,32'd1969344934,32'd2534523080,32'd2665563904,32'd3514892628,32'd265049099,32'd2449404120,32'd453065119,32'd3795864463,32'd1569683418,32'd539639323,32'd2287008439,32'd3972660041,32'd1730605673,32'd480498390,32'd1007512487,32'd3318166191,32'd3796449494,32'd3449856475,32'd1717914918,32'd2795959904,32'd45383166,32'd485558549,32'd3950876764,32'd1634068959,32'd896867387,32'd1917283619,32'd3953675561,32'd1187332833,32'd1994019922,32'd4268194620,32'd4102008957,32'd936120505,32'd1294478167,32'd3841025952,32'd1699618892,32'd2194081082,32'd611750005,32'd2147383559,32'd2231395445,32'd1983126147,32'd2265109737,32'd141910303,32'd161423763,32'd462233764,32'd2632116865,32'd3757086488,32'd4212233956,32'd1125914118,32'd3660165513,32'd3457529378,32'd2732673041,32'd860032883,32'd2064802063,32'd3799566677,32'd843058885,32'd597068400,32'd3542060425,32'd359920673,32'd4110743408,32'd4050317728,32'd1892992132,32'd2934259476,32'd1550715292,32'd1706316388,32'd3109212504,32'd954907921,32'd3825832114,32'd1854233928,32'd4001025594,32'd1406585576,32'd3968201444,32'd2577977181,32'd2655923113,32'd3421075971,32'd1088809168,32'd3881027887,32'd1051168756,32'd2986286440,32'd981744121,32'd3569720512,32'd313287791,32'd2575857120,32'd1301784708,32'd314202987,32'd3132941411,32'd1240723705,32'd1391137252,32'd2671656400,32'd325625733,32'd3696778854,32'd284461833,32'd3202770816,32'd3941535311,32'd607643288,32'd2529629289,32'd1371755819,32'd1489632964,32'd1012800992,32'd2670621135,32'd1832011890,32'd281952627,32'd610765913,32'd3925701436,32'd106823192,32'd4226412442,32'd282321962,32'd3215726425,32'd3356372094,32'd2328724316,32'd127157074,32'd2230415839,32'd2932373212,32'd3590303986,32'd4227905160,32'd767063856,32'd614167064,32'd1605707990,32'd1975939317,32'd2771236582,32'd1137581788,32'd980888698,32'd2808583945,32'd2266356233,32'd3714884555,32'd3683686884,32'd3562644229,32'd2462549847,32'd3775753525,32'd2844284824,32'd1958640221,32'd2354026721,32'd2054107185,32'd3264939860,32'd1112874779,32'd3956938481,32'd2037033584,32'd2280810156,32'd2067589016,32'd2603507610,32'd1175446314,32'd2718629137,32'd698822522,32'd2224934154,32'd2297021184,32'd2693039652,32'd3780746374,32'd3614057572,32'd367436315,32'd3763313683,32'd3505045078,32'd2831416447,32'd3535515583,32'd4277891831,32'd837664826,32'd3932714317,32'd961491174,32'd2127070362,32'd2693520819,32'd198269976,32'd1311855742,32'd3566819907,32'd2347785709,32'd2566048980,32'd3557034492,32'd2783662465,32'd676528503,32'd2373484829,32'd840509954,32'd3519123538,32'd2625414289,32'd1566383306,32'd836340051,32'd2478087736,32'd2840453856,32'd1855512191,32'd95009460,32'd1555072155,32'd1030225246,32'd2877123406,32'd94227745,32'd2882166470,32'd3806317775,32'd1926821318,32'd2250056281,32'd3382188205,32'd4088822114,32'd1223816410,32'd3072671496,32'd1613109469,32'd2143978386,32'd4009374062,32'd262993567,32'd2753953039,32'd1300608482,32'd2385138085,32'd1233652508,32'd1220770796,32'd1476834675,32'd102614847,32'd3870616539,32'd2935588114,32'd1653162115,32'd2818865106,32'd3576835843,32'd4213508374,32'd3434980330,32'd1720449988,32'd4033654965,32'd3740957436,32'd2386309702,32'd3539167101,32'd1140754642,32'd4123661669,32'd1392372379,32'd376204646,32'd3898673786,32'd1886893516,32'd2891199990,32'd437801529,32'd2923086221,32'd3810238677,32'd2449469876,32'd1479383443,32'd2814550949,32'd2440339870,32'd3131865469,32'd732815996,32'd1036426282,32'd597866774,32'd2216566078,32'd607322300,32'd4050607484,32'd1454330362,32'd3155158821,32'd1638923698,32'd179684232,32'd2536571847,32'd2413832827,32'd1581410039,32'd2164382601,32'd2292163827,32'd3746505897,32'd3096953148,32'd2640545275,32'd3286135343,32'd3191454495,32'd3228651068,32'd3588672187,32'd3452239013,32'd1592291796,32'd2973452884,32'd1812273278,32'd1709930435,32'd3661313599,32'd4224925813,32'd3540177092,32'd2002781766,32'd4201769589,32'd2676817993,32'd1349669984,32'd2906395199,32'd4019597455,32'd1345782310,32'd921967201,32'd2598854474,32'd2667646161,32'd1948434636,32'd3784365245,32'd1145213362,32'd3224868746,32'd2402025379,32'd3364128315,32'd1785085746,32'd92883131,32'd3306961981,32'd792772838,32'd4033622241,32'd681580311,32'd2983301384,32'd2629073562};
end
else begin
	if(enable)out<=in;
end
endmodule